
// === Extension board configuration ===
// Uncomment the following define if you have the HX8K Breakout Board Extension.
// Information about that extension board:
//    https://github.com/maikmerten/hx8k-breakout-extension
// With the extension board present, RAM capacity is 512 KB.
// Without the extension board, RAM capacity is 8 KB.

`define EXTENSION_PRESENT

